magic
tech sky130A
magscale 1 2
timestamp 1647132523
<< nwell >>
rect 228 -171 546 316
<< pwell >>
rect -294 -170 228 316
<< nmos >>
rect -160 186 160 216
rect -160 100 160 130
<< pmos >>
rect 264 186 510 216
rect 264 100 510 130
<< ndiff >>
rect -160 261 160 269
rect -160 227 -117 261
rect -83 227 -49 261
rect -15 227 19 261
rect 53 227 87 261
rect 121 227 160 261
rect -160 216 160 227
rect -160 130 160 186
rect -160 89 160 100
rect -160 55 -119 89
rect -85 55 -51 89
rect -17 55 17 89
rect 51 55 85 89
rect 119 55 160 89
rect -160 47 160 55
<< pdiff >>
rect 264 261 510 269
rect 264 227 302 261
rect 336 227 370 261
rect 404 227 438 261
rect 472 227 510 261
rect 264 216 510 227
rect 264 175 510 186
rect 264 141 302 175
rect 336 141 370 175
rect 404 141 438 175
rect 472 141 510 175
rect 264 130 510 141
rect 264 89 510 100
rect 264 55 302 89
rect 336 55 370 89
rect 404 55 438 89
rect 472 55 510 89
rect 264 47 510 55
<< ndiffc >>
rect -117 227 -83 261
rect -49 227 -15 261
rect 19 227 53 261
rect 87 227 121 261
rect -119 55 -85 89
rect -51 55 -17 89
rect 17 55 51 89
rect 85 55 119 89
<< pdiffc >>
rect 302 227 336 261
rect 370 227 404 261
rect 438 227 472 261
rect 302 141 336 175
rect 370 141 404 175
rect 438 141 472 175
rect 302 55 336 89
rect 370 55 404 89
rect 438 55 472 89
<< psubdiff >>
rect -95 -67 76 -54
rect -95 -101 -20 -67
rect 14 -101 76 -67
rect -95 -114 76 -101
<< nsubdiff >>
rect 319 -21 452 -10
rect 319 -55 368 -21
rect 402 -55 452 -21
rect 319 -77 452 -55
<< psubdiffcont >>
rect -20 -101 14 -67
<< nsubdiffcont >>
rect 368 -55 402 -21
<< poly >>
rect -252 230 -186 240
rect -252 196 -236 230
rect -202 216 -186 230
rect -202 196 -160 216
rect -252 186 -160 196
rect 160 186 264 216
rect 510 186 536 216
rect -252 120 -160 130
rect -252 86 -236 120
rect -202 100 -160 120
rect 160 100 264 130
rect 510 100 536 130
rect -202 86 -186 100
rect -252 76 -186 86
<< polycont >>
rect -236 196 -202 230
rect -236 86 -202 120
<< locali >>
rect -236 230 -202 246
rect -160 227 -117 261
rect -83 227 -49 261
rect -15 227 19 261
rect 53 227 87 261
rect 121 227 302 261
rect 336 227 370 261
rect 404 227 438 261
rect 472 227 546 261
rect -236 180 -202 196
rect -236 120 -202 136
rect 195 89 229 227
rect 264 141 302 175
rect 336 141 370 175
rect 404 141 438 175
rect 472 141 510 175
rect -236 70 -202 86
rect -160 55 -119 89
rect -85 55 -51 89
rect 51 55 85 89
rect 119 55 160 89
rect 195 55 302 89
rect 336 55 370 89
rect 404 55 438 89
rect 472 55 546 89
rect 346 -21 431 -11
rect -95 -67 76 -54
rect 346 -55 368 -21
rect 402 -55 431 -21
rect 346 -64 431 -55
rect -95 -101 -20 -67
rect 14 -101 76 -67
rect -95 -114 76 -101
<< viali >>
rect 370 141 404 175
rect -17 55 17 89
rect 368 -55 402 -21
rect -20 -101 14 -67
<< metal1 >>
rect -29 89 29 316
rect -29 55 -17 89
rect 17 55 29 89
rect -29 -67 29 55
rect -29 -101 -20 -67
rect 14 -101 29 -67
rect -29 -144 29 -101
rect 358 175 416 316
rect 358 141 370 175
rect 404 141 416 175
rect 358 -21 416 141
rect 358 -55 368 -21
rect 402 -55 416 -21
rect 358 -112 416 -55
<< labels >>
rlabel locali -236 70 -202 136 7 B
port 1 w
rlabel locali -236 180 -202 246 7 A
port 0 w
rlabel locali -160 227 546 261 3 Y
port 4 e
rlabel metal1 -29 0 29 316 5 VGND
port 2 s
rlabel metal1 358 0 416 316 1 VPWR
port 3 n
rlabel nwell 228 0 546 316 3 VPB
<< end >>
